library ieee;

use ieee.std_logic_1164.all;
use.ieee.std.logic_unsigned.all;

entity decoder is

    port   (
            -- clock : in std_logic;
            dataOut : std_logic_vector ( 31 down to 0);
            instruction : out std_logic_vector ( 4 down to 0);
            immediat : out std_logic_vector ( 15 down to 0);
            operator1 : out std_logic_vector ( 7 down to 0);
            operator2 : out std_logic_vector ( 7 down to 0);
            operator3 : out std_logic_vector ( 7 down to 0);
            )

end entity decoder;

architecture decode of decoder is


    begin

        instruction <= dataOut(31 to 27);

        if (instructuin = 1)
            then
                if dataOut(26) = x"1" ....
                else ...

        elseif (instructuin = x)
            then
                if dataOut(26) = x"1" ....
                else ...

        elseif(instructuin=2)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=3)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=4)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=5)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=6)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=7)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=8)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=9)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=10)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=11)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=12)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=13)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=14)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=15)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=16)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=17)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif(instructuin=18)
            then
                if dataOut(26) = x"1"....
                else ...

        elseif

-- elseif(instructuin=XXXXX)
-- then
-- if dataOut(26) = x"1"....
-- else ...

    end

end architecture decode;
