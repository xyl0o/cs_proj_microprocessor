package constants is
	constant data_len: integer := 32;
end package constants;