package constants is
	constant data_len: integer := 32;
	constant immediate_len: integer := 16;
	constant reg_addr_len: integer := 6;
	constant op_code_len: integer := 5;
	constant alu_op_code_len: integer := 5;
end package constants;