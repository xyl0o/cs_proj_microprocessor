regType is array (0 to 31) of std_logic_vector(31 downto 0);

